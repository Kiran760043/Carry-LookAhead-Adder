//////////////////////////////////////////////////////////////////////////////////
// Design Name: Full Adder for GP
// Engineer: kiran
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps


module full_adder_gp(
    input  wire A,
    input  wire B,
    input  wire Ci,
    output wire S,
    output wire Co
    );

    assign S  = A ^ B ^ Ci;

endmodule
